//`define NEW_19811_USB_CORES

`ifndef NEW_19811_USB_CORES
module usb_gowin_top (
    input  wire        clk480_i      ,
    input  wire        clk60_i       ,
    input  wire        rst_i         ,
    input  wire        pll_lock_i    ,

    usb_gowin_if.gwn   usb            ,
    output wire        utmi_txvalid_o ,
    output wire        utmi_txready_o ,

    inout  wire        usb_dxp_io      ,
    inout  wire        usb_dxn_io      ,
    input  wire        usb_rxdp_i      ,
    input  wire        usb_rxdn_i      ,
    output wire        usb_pullup_en_o ,
    inout  wire        usb_term_dp_io  ,
    inout  wire        usb_term_dn_io
    ,output wire w_eop_o
    ,output wire [3:0]  q_offset_o 
    ,output wire [3:0] crc_dbg_dataout_o
    ,output wire stuck_in_2nd_or_3rd_state_o
    ,output wire [15 : 0] DRU_dbg_signals_o
    ,output wire [19 : 0] dev_controller_dbg_o
);

    wire [1:0]  PHY_XCVRSELECT;
    wire        PHY_TERMSELECT;
    wire [1:0]  PHY_OPMODE;
    wire [1:0]  PHY_LINESTATE;
    wire        PHY_TXVALID;
    wire        PHY_TXREADY;
    wire        PHY_RXVALID;
    wire        PHY_RXACTIVE;
    wire        PHY_RXERROR;
    wire [7:0]  PHY_DATAIN;
    wire [7:0]  PHY_DATAOUT;
    wire        PHY_RESET;

    wire [9:0]  DESCROM_RADDR;
    wire [7:0]  DESCROM_RDAT;
    wire [9:0]  DESC_DEV_ADDR;
    wire [7:0]  DESC_DEV_LEN;
    wire [9:0]  DESC_QUAL_ADDR;
    wire [7:0]  DESC_QUAL_LEN;
    wire [9:0]  DESC_FSCFG_ADDR;
    wire [7:0]  DESC_FSCFG_LEN;
    wire [9:0]  DESC_HSCFG_ADDR;
    wire [7:0]  DESC_HSCFG_LEN;
    wire [9:0]  DESC_OSCFG_ADDR;
    wire [9:0]  DESC_STRLANG_ADDR;
    wire [9:0]  DESC_STRVENDOR_ADDR;
    wire [7:0]  DESC_STRVENDOR_LEN;
    wire [9:0]  DESC_STRPRODUCT_ADDR;
    wire [7:0]  DESC_STRPRODUCT_LEN;
    wire [9:0]  DESC_STRSERIAL_ADDR;
    wire [7:0]  DESC_STRSERIAL_LEN;
    wire        DESCROM_HAVE_STRINGS;
    wire sclk;

    USB_Device_Controller_Top u_usb_device_controller_top (
        .clk_i                 ( clk60_i             ),
        .reset_i               ( rst_i                ),
        .usbrst_o              (                        ),
        .highspeed_o           (                        ),
        .suspend_o             (                        ),
        .online_o              (                        ),
        .txdat_i               ( usb.txdat ),
        .txval_i               ( usb.txval ),
        .txdat_len_i           ( usb.txdat_len ),
        .txcork_i              ( usb.txcork ),
        .txiso_pid_i           ( 4'b0000                ),
        .txpop_o               ( usb.txpop ),
        .txact_o               ( usb.txact ),
        .txpktfin_o            (                        ),
        .rxdat_o               ( usb.rxdat ),
        .rxval_o               ( usb.rxval ),
        .rxact_o               ( usb.rxact ),
        .rxrdy_i               ( usb.rxrdy ),
        .rxpktval_o            (                        ),
        .setup_o               ( usb.setup ),
        .endpt_o               ( usb.endpt ),
        .sof_o                 (                        ),
        .inf_alter_i           ( 8'd0                   ),
        .inf_alter_o           (                        ),
        .inf_sel_o             (                        ),
        .inf_set_o             (                        ),
        .descrom_rdata_i       ( DESCROM_RDAT           ),
        .descrom_raddr_o       ( DESCROM_RADDR          ),
        .desc_dev_addr_i       ( DESC_DEV_ADDR          ),
        .desc_dev_len_i        ( DESC_DEV_LEN           ),
        .desc_qual_addr_i      ( DESC_QUAL_ADDR         ),
        .desc_qual_len_i       ( DESC_QUAL_LEN          ),
        .desc_fscfg_addr_i     ( DESC_FSCFG_ADDR        ),
        .desc_fscfg_len_i      ( DESC_FSCFG_LEN         ),
        .desc_hscfg_addr_i     ( DESC_HSCFG_ADDR        ),
        .desc_hscfg_len_i      ( DESC_HSCFG_LEN         ),
        .desc_oscfg_addr_i     ( DESC_OSCFG_ADDR        ),
        .desc_strlang_addr_i   ( DESC_STRLANG_ADDR      ),
        .desc_strvendor_addr_i ( DESC_STRVENDOR_ADDR    ),
        .desc_strvendor_len_i  ( DESC_STRVENDOR_LEN     ),
        .desc_strproduct_addr_i( DESC_STRPRODUCT_ADDR   ),
        .desc_strproduct_len_i ( DESC_STRPRODUCT_LEN    ),
        .desc_strserial_addr_i ( DESC_STRSERIAL_ADDR    ),
        .desc_strserial_len_i  ( DESC_STRSERIAL_LEN     ),
        .desc_have_strings_i   ( DESCROM_HAVE_STRINGS   ),
        .utmi_dataout_o        ( PHY_DATAOUT            ),
        .utmi_txvalid_o        ( PHY_TXVALID            ),
        .utmi_txready_i        ( PHY_TXREADY            ),
        .utmi_datain_i         ( PHY_DATAIN             ),
        .utmi_rxactive_i       ( PHY_RXACTIVE           ),
        .utmi_rxvalid_i        ( PHY_RXVALID            ),
        .utmi_rxerror_i        ( PHY_RXERROR            ),
        .utmi_linestate_i      ( PHY_LINESTATE          ),
        .utmi_opmode_o         ( PHY_OPMODE             ),
        .utmi_xcvrselect_o     ( PHY_XCVRSELECT         ),
        .utmi_termselect_o     ( PHY_TERMSELECT         ),
        .utmi_reset_o          ( PHY_RESET              ),
        .ack_timeout_o         ( usb.ack_tout           ),
        .ack_received_o        ( usb.ack_received       ),
        .ack_bad_packet_o      ( usb.ack_bad_packet     )
        ,.transact_state_o (usb.transact_state_o)
        ,.clk_120              ( sclk)
        ,.crc_dbg_dataout_o (crc_dbg_dataout_o)
        ,.stuck_in_2nd_or_3rd_state_o (stuck_in_2nd_or_3rd_state_o)
        ,.dev_controller_dbg_o        (dev_controller_dbg_o)
    );

`ifdef USB_CDC_ENA
    usb_desc_msd_cdc #(
        .VENDORID    ( 16'h33AA ),
        .PRODUCTID   ( 16'h0000 ),
        .VERSIONBCD  ( 16'h0100 ),
        .HSSUPPORT   ( 1        ),
        .SELFPOWERED ( 1        )
    ) u_usb_desc (
            .CLK                    ( clk60_i           ) ,
            .RESET                  ( rst_i              ) ,
            .i_pid                  ( 16'd0                ) ,
            .i_vid                  ( 16'd0                ) ,
            .i_descrom_raddr        ( DESCROM_RADDR        ) ,
            .o_descrom_rdat         ( DESCROM_RDAT         ) ,
            .o_desc_dev_addr        ( DESC_DEV_ADDR        ) ,
            .o_desc_dev_len         ( DESC_DEV_LEN         ) ,
            .o_desc_qual_addr       ( DESC_QUAL_ADDR       ) ,
            .o_desc_qual_len        ( DESC_QUAL_LEN        ) ,
            .o_desc_fscfg_addr      ( DESC_FSCFG_ADDR      ) ,
            .o_desc_fscfg_len       ( DESC_FSCFG_LEN       ) ,
            .o_desc_hscfg_addr      ( DESC_HSCFG_ADDR      ) ,
            .o_desc_hscfg_len       ( DESC_HSCFG_LEN       ) ,
            .o_desc_oscfg_addr      ( DESC_OSCFG_ADDR      ) ,
            .o_desc_strlang_addr    ( DESC_STRLANG_ADDR    ) ,
            .o_desc_strvendor_addr  ( DESC_STRVENDOR_ADDR  ) ,
            .o_desc_strvendor_len   ( DESC_STRVENDOR_LEN   ) ,
            .o_desc_strproduct_addr ( DESC_STRPRODUCT_ADDR ) ,
            .o_desc_strproduct_len  ( DESC_STRPRODUCT_LEN  ) ,
            .o_desc_strserial_addr  ( DESC_STRSERIAL_ADDR  ) ,
            .o_desc_strserial_len   ( DESC_STRSERIAL_LEN   ) ,
            .o_descrom_have_strings ( DESCROM_HAVE_STRINGS )
    );
`else
    usb_desc_msd #(
        .VENDORID    ( 16'h33AA ),
        .PRODUCTID   ( 16'h0000 ),
        .VERSIONBCD  ( 16'h0100 ),
        .HSSUPPORT   ( 1        ),
        .SELFPOWERED ( 1        )
    ) u_usb_desc (
            .CLK                    ( clk60_i           ) ,
            .RESET                  ( rst_i              ) ,
            .i_pid                  ( 16'd0                ) ,
            .i_vid                  ( 16'd0                ) ,
            .i_descrom_raddr        ( DESCROM_RADDR        ) ,
            .o_descrom_rdat         ( DESCROM_RDAT         ) ,
            .o_desc_dev_addr        ( DESC_DEV_ADDR        ) ,
            .o_desc_dev_len         ( DESC_DEV_LEN         ) ,
            .o_desc_qual_addr       ( DESC_QUAL_ADDR       ) ,
            .o_desc_qual_len        ( DESC_QUAL_LEN        ) ,
            .o_desc_fscfg_addr      ( DESC_FSCFG_ADDR      ) ,
            .o_desc_fscfg_len       ( DESC_FSCFG_LEN       ) ,
            .o_desc_hscfg_addr      ( DESC_HSCFG_ADDR      ) ,
            .o_desc_hscfg_len       ( DESC_HSCFG_LEN       ) ,
            .o_desc_oscfg_addr      ( DESC_OSCFG_ADDR      ) ,
            .o_desc_strlang_addr    ( DESC_STRLANG_ADDR    ) ,
            .o_desc_strvendor_addr  ( DESC_STRVENDOR_ADDR  ) ,
            .o_desc_strvendor_len   ( DESC_STRVENDOR_LEN   ) ,
            .o_desc_strproduct_addr ( DESC_STRPRODUCT_ADDR ) ,
            .o_desc_strproduct_len  ( DESC_STRPRODUCT_LEN  ) ,
            .o_desc_strserial_addr  ( DESC_STRSERIAL_ADDR  ) ,
            .o_desc_strserial_len   ( DESC_STRSERIAL_LEN   ) ,
            .o_descrom_have_strings ( DESCROM_HAVE_STRINGS )
    );
`endif

    USB2_0_SoftPHY_Top u_USB_SoftPHY_Top (
        .clk_i            (clk60_i     ),
        .rst_i            (PHY_RESET      ),
        .fclk_i           (clk480_i    ),
        .pll_locked_i     (pll_lock_i     ),

        .utmi_data_out_i  (PHY_DATAOUT    ),
        .utmi_txvalid_i   (PHY_TXVALID    ),
        .utmi_op_mode_i   (PHY_OPMODE     ),
        .utmi_xcvrselect_i(PHY_XCVRSELECT ),
        .utmi_termselect_i(PHY_TERMSELECT ),
        .utmi_data_in_o   (PHY_DATAIN     ),
        .utmi_txready_o   (PHY_TXREADY    ),
        .utmi_rxvalid_o   (PHY_RXVALID    ),
        .utmi_rxactive_o  (PHY_RXACTIVE   ),
        .utmi_rxerror_o   (PHY_RXERROR    ),
        .utmi_linestate_o (PHY_LINESTATE  ),

        .usb_dxp_io       (usb_dxp_io     ),
        .usb_dxn_io       (usb_dxn_io     ),
        .usb_rxdp_i       (usb_rxdp_i     ),
        .usb_rxdn_i       (usb_rxdn_i     ),
        .usb_pullup_en_o  (usb_pullup_en_o),
        .usb_term_dp_io   (usb_term_dp_io ),
        .usb_term_dn_io   (usb_term_dn_io )
        ,.w_eop_o         (w_eop_o)
        ,.q_offset_o      (q_offset_o)
        ,.sclk            (sclk)
        ,.DRU_dbg_signals_o(DRU_dbg_signals_o)
    );

    assign utmi_txvalid_o = PHY_TXVALID ;
    assign utmi_txready_o = PHY_TXREADY ;
endmodule










`else


















module usb_gowin_top (
    input  wire        clk480_i      ,
    input  wire        clk60_i       ,
    input  wire        rst_i         ,
    input  wire        pll_lock_i    ,

    usb_gowin_if.gwn   usb            ,
    output wire        utmi_txvalid_o ,
    output wire        utmi_txready_o ,

    inout  wire        usb_dxp_io      ,
    inout  wire        usb_dxn_io      ,
    input  wire        usb_rxdp_i      ,
    input  wire        usb_rxdn_i      ,
    output wire        usb_pullup_en_o ,
    inout  wire        usb_term_dp_io  ,
    inout  wire        usb_term_dn_io
    ,output wire w_eop_o
    ,output wire [3:0]  q_offset_o 
    ,output wire [3:0] crc_dbg_dataout_o
    ,output wire stuck_in_2nd_or_3rd_state_o
    ,output wire [15 : 0] DRU_dbg_signals_o
    ,output wire [19 : 0] dev_controller_dbg_o
);

    wire [1:0]  PHY_XCVRSELECT;
    wire        PHY_TERMSELECT;
    wire [1:0]  PHY_OPMODE;
    wire [1:0]  PHY_LINESTATE;
    wire        PHY_TXVALID;
    wire        PHY_TXREADY;
    wire        PHY_RXVALID;
    wire        PHY_RXACTIVE;
    wire        PHY_RXERROR;
    wire [7:0]  PHY_DATAIN;
    wire [7:0]  PHY_DATAOUT;
    wire        PHY_RESET;

    wire [9:0]  DESCROM_RADDR;
    wire [7:0]  DESCROM_RDAT;
    wire [9:0]  DESC_DEV_ADDR;
    wire [7:0]  DESC_DEV_LEN;
    wire [9:0]  DESC_QUAL_ADDR;
    wire [7:0]  DESC_QUAL_LEN;
    wire [9:0]  DESC_FSCFG_ADDR;
    wire [7:0]  DESC_FSCFG_LEN;
    wire [9:0]  DESC_HSCFG_ADDR;
    wire [7:0]  DESC_HSCFG_LEN;
    wire [9:0]  DESC_OSCFG_ADDR;
    wire [9:0]  DESC_STRLANG_ADDR;
    wire [9:0]  DESC_STRVENDOR_ADDR;
    wire [7:0]  DESC_STRVENDOR_LEN;
    wire [9:0]  DESC_STRPRODUCT_ADDR;
    wire [7:0]  DESC_STRPRODUCT_LEN;
    wire [9:0]  DESC_STRSERIAL_ADDR;
    wire [7:0]  DESC_STRSERIAL_LEN;
    wire        DESCROM_HAVE_STRINGS;
    wire sclk;

    USB_Device_Controller_Top u_usb_device_controller_top (
        .clk_i                 ( clk60_i             ),
        .reset_i               ( rst_i                ),
        .usbrst_o              (                        ),
        .highspeed_o           (                        ),
        .suspend_o             (                        ),
        .online_o              (                        ),
        .txdat_i               ( usb.txdat ),
        .txval_i               ( usb.txval ),
        .txdat_len_i           ( usb.txdat_len ),
        .txcork_i              ( usb.txcork ),
        .txiso_pid_i           ( 4'b0000                ),
        .txpop_o               ( usb.txpop ),
        .txact_o               ( usb.txact ),
        .txpktfin_o            (                        ),
        .rxdat_o               ( usb.rxdat ),
        .rxval_o               ( usb.rxval ),
        .rxact_o               ( usb.rxact ),
        .rxrdy_i               ( usb.rxrdy ),
        .rxpktval_o            (                        ),
        .setup_o               ( usb.setup ),
        .endpt_o               ( usb.endpt ),
        .sof_o                 (                        ),
        .inf_alter_i           ( 8'd0                   ),
        .inf_alter_o           (                        ),
        .inf_sel_o             (                        ),
        .inf_set_o             (                        ),
        .descrom_rdata_i       ( DESCROM_RDAT           ),
        .descrom_raddr_o       ( DESCROM_RADDR          ),
        .desc_dev_addr_i       ( DESC_DEV_ADDR          ),
        .desc_dev_len_i        ( DESC_DEV_LEN           ),
        .desc_qual_addr_i      ( DESC_QUAL_ADDR         ),
        .desc_qual_len_i       ( DESC_QUAL_LEN          ),
        .desc_fscfg_addr_i     ( DESC_FSCFG_ADDR        ),
        .desc_fscfg_len_i      ( DESC_FSCFG_LEN         ),
        .desc_hscfg_addr_i     ( DESC_HSCFG_ADDR        ),
        .desc_hscfg_len_i      ( DESC_HSCFG_LEN         ),
        .desc_oscfg_addr_i     ( DESC_OSCFG_ADDR        ),
        .desc_strlang_addr_i   ( DESC_STRLANG_ADDR      ),
        .desc_strvendor_addr_i ( DESC_STRVENDOR_ADDR    ),
        .desc_strvendor_len_i  ( DESC_STRVENDOR_LEN     ),
        .desc_strproduct_addr_i( DESC_STRPRODUCT_ADDR   ),
        .desc_strproduct_len_i ( DESC_STRPRODUCT_LEN    ),
        .desc_strserial_addr_i ( DESC_STRSERIAL_ADDR    ),
        .desc_strserial_len_i  ( DESC_STRSERIAL_LEN     ),
        .desc_have_strings_i   ( DESCROM_HAVE_STRINGS   ),
        .utmi_dataout_o        ( PHY_DATAOUT            ),
        .utmi_txvalid_o        ( PHY_TXVALID            ),
        .utmi_txready_i        ( PHY_TXREADY            ),
        .utmi_datain_i         ( PHY_DATAIN             ),
        .utmi_rxactive_i       ( PHY_RXACTIVE           ),
        .utmi_rxvalid_i        ( PHY_RXVALID            ),
        .utmi_rxerror_i        ( PHY_RXERROR            ),
        .utmi_linestate_i      ( PHY_LINESTATE          ),
        .utmi_opmode_o         ( PHY_OPMODE             ),
        .utmi_xcvrselect_o     ( PHY_XCVRSELECT         ),
        .utmi_termselect_o     ( PHY_TERMSELECT         ),
        .utmi_reset_o          ( PHY_RESET              )
    );

`ifdef USB_CDC_ENA
    usb_desc_msd_cdc #(
        .VENDORID    ( 16'h33AA ),
        .PRODUCTID   ( 16'h0000 ),
        .VERSIONBCD  ( 16'h0100 ),
        .HSSUPPORT   ( 1        ),
        .SELFPOWERED ( 1        )
    ) u_usb_desc (
            .CLK                    ( clk60_i           ) ,
            .RESET                  ( rst_i              ) ,
            .i_pid                  ( 16'd0                ) ,
            .i_vid                  ( 16'd0                ) ,
            .i_descrom_raddr        ( DESCROM_RADDR        ) ,
            .o_descrom_rdat         ( DESCROM_RDAT         ) ,
            .o_desc_dev_addr        ( DESC_DEV_ADDR        ) ,
            .o_desc_dev_len         ( DESC_DEV_LEN         ) ,
            .o_desc_qual_addr       ( DESC_QUAL_ADDR       ) ,
            .o_desc_qual_len        ( DESC_QUAL_LEN        ) ,
            .o_desc_fscfg_addr      ( DESC_FSCFG_ADDR      ) ,
            .o_desc_fscfg_len       ( DESC_FSCFG_LEN       ) ,
            .o_desc_hscfg_addr      ( DESC_HSCFG_ADDR      ) ,
            .o_desc_hscfg_len       ( DESC_HSCFG_LEN       ) ,
            .o_desc_oscfg_addr      ( DESC_OSCFG_ADDR      ) ,
            .o_desc_strlang_addr    ( DESC_STRLANG_ADDR    ) ,
            .o_desc_strvendor_addr  ( DESC_STRVENDOR_ADDR  ) ,
            .o_desc_strvendor_len   ( DESC_STRVENDOR_LEN   ) ,
            .o_desc_strproduct_addr ( DESC_STRPRODUCT_ADDR ) ,
            .o_desc_strproduct_len  ( DESC_STRPRODUCT_LEN  ) ,
            .o_desc_strserial_addr  ( DESC_STRSERIAL_ADDR  ) ,
            .o_desc_strserial_len   ( DESC_STRSERIAL_LEN   ) ,
            .o_descrom_have_strings ( DESCROM_HAVE_STRINGS )
    );
`else
    usb_desc_msd #(
        .VENDORID    ( 16'h33AA ),
        .PRODUCTID   ( 16'h0000 ),
        .VERSIONBCD  ( 16'h0100 ),
        .HSSUPPORT   ( 1        ),
        .SELFPOWERED ( 1        )
    ) u_usb_desc (
            .CLK                    ( clk60_i           ) ,
            .RESET                  ( rst_i              ) ,
            .i_pid                  ( 16'd0                ) ,
            .i_vid                  ( 16'd0                ) ,
            .i_descrom_raddr        ( DESCROM_RADDR        ) ,
            .o_descrom_rdat         ( DESCROM_RDAT         ) ,
            .o_desc_dev_addr        ( DESC_DEV_ADDR        ) ,
            .o_desc_dev_len         ( DESC_DEV_LEN         ) ,
            .o_desc_qual_addr       ( DESC_QUAL_ADDR       ) ,
            .o_desc_qual_len        ( DESC_QUAL_LEN        ) ,
            .o_desc_fscfg_addr      ( DESC_FSCFG_ADDR      ) ,
            .o_desc_fscfg_len       ( DESC_FSCFG_LEN       ) ,
            .o_desc_hscfg_addr      ( DESC_HSCFG_ADDR      ) ,
            .o_desc_hscfg_len       ( DESC_HSCFG_LEN       ) ,
            .o_desc_oscfg_addr      ( DESC_OSCFG_ADDR      ) ,
            .o_desc_strlang_addr    ( DESC_STRLANG_ADDR    ) ,
            .o_desc_strvendor_addr  ( DESC_STRVENDOR_ADDR  ) ,
            .o_desc_strvendor_len   ( DESC_STRVENDOR_LEN   ) ,
            .o_desc_strproduct_addr ( DESC_STRPRODUCT_ADDR ) ,
            .o_desc_strproduct_len  ( DESC_STRPRODUCT_LEN  ) ,
            .o_desc_strserial_addr  ( DESC_STRSERIAL_ADDR  ) ,
            .o_desc_strserial_len   ( DESC_STRSERIAL_LEN   ) ,
            .o_descrom_have_strings ( DESCROM_HAVE_STRINGS )
    );
`endif

    USB2_0_SoftPHY_Top u_USB_SoftPHY_Top (
        .clk_i            (clk60_i     ),
        .rst_i            (PHY_RESET      ),
        .fclk_i           (clk480_i    ),
        .pll_locked_i     (pll_lock_i     ),

        .utmi_data_out_i  (PHY_DATAOUT    ),
        .utmi_txvalid_i   (PHY_TXVALID    ),
        .utmi_op_mode_i   (PHY_OPMODE     ),
        .utmi_xcvrselect_i(PHY_XCVRSELECT ),
        .utmi_termselect_i(PHY_TERMSELECT ),
        .utmi_data_in_o   (PHY_DATAIN     ),
        .utmi_txready_o   (PHY_TXREADY    ),
        .utmi_rxvalid_o   (PHY_RXVALID    ),
        .utmi_rxactive_o  (PHY_RXACTIVE   ),
        .utmi_rxerror_o   (PHY_RXERROR    ),
        .utmi_linestate_o (PHY_LINESTATE  ),

        .usb_dxp_io       (usb_dxp_io     ),
        .usb_dxn_io       (usb_dxn_io     ),
        .usb_rxdp_i       (usb_rxdp_i     ),
        .usb_rxdn_i       (usb_rxdn_i     ),
        .usb_pullup_en_o  (usb_pullup_en_o),
        .usb_term_dp_io   (usb_term_dp_io ),
        .usb_term_dn_io   (usb_term_dn_io )
    );

    assign utmi_txvalid_o = PHY_TXVALID ;
    assign utmi_txready_o = PHY_TXREADY ;
endmodule
`endif
